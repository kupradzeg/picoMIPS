//-----------------------------------------------------	
//	File	Name			:	alucodes.sv	
//	FuncRon				:	pMIPS	ALU	funcRon	code	definiRons		
//	Author:			tjk
//	Last	rev.	23	Oct	12		
//-----------------------------------------------------	
//		
`define	RA			2'b00	
`define	RB			2'b01	
`define	RADD		2'b10	
`define	RMUL		2'b11			
