//-----------------------------------------------------
// File Name   : alu.sv
// Function    : ALU module for picoMIPS
// Version: 1,  only 8 funcs
// Author:  tjk
// Last rev. 23 Oct 12
//-----------------------------------------------------

`include "alucodes.sv"  
//`include "mult.sv"
module alu #(parameter n =8) (
   input logic signed [n-1:0] a, b, // ALU operands
   input logic [1:0] func, // ALU function code

   output logic signed [n-1:0] result // ALU result
);       
//------------- code starts here ---------
 
// Instantiate the multiplier module
logic signed [n*2-1:0] temp;
signed_mult multiplier(.out(temp), .a(a), .b(b));
 
// create the ALU, use signal ar in arithmetic operations
always_comb
begin
  //default output values; prevent latches 

  result = a; // default
   
  case(func)
  	`RA   : result = a;
	`RB   : result = b;
     `RADD  : begin
	     result = a+b; // arithmetic addition

		end
	`RMUL: begin
		
		result = temp[14:7];
	end

   endcase
	 
 
 
 end //always_comb

endmodule //end of module ALU


