//-----------------------------------------------------	
//	File	Name			:	opcodes.sv	
//	FuncRon				:	pMIPS	ALU	funcRon	code	definiRons		
//	Author:			tjk
//	Last	rev.	23	Oct	12		
//-----------------------------------------------------	
//		

`define ST_0	5'b00000
`define ST_1	5'b00100
`define ADD		5'b01010 
`define ADDI	5'b01110
`define MUL		5'b10011
`define MULI	5'b10111
`define	IMM		5'b11001 
`define SWI		5'b11101